module cond_sub
	(
		input wire[3:0] i,
		output wire [3:0] o
	);
	
	assign o =
				(i == 4'b0000) ? 4'b0000 :
				(i == 4'b0001) ? 4'b0001 :
				(i == 4'b0010) ? 4'b0010 :
				(i == 4'b0011) ? 4'b0011 :
				(i == 4'b0100) ? 4'b0100 :
				(i == 4'b1000) ? 4'b0101 :
				(i == 4'b1001) ? 4'b0110 :
				(i == 4'b1010) ? 4'b0111 :
				(i == 4'b1011) ? 4'b1000 :
				(i == 4'b1100) ? 4'b1001 :
									  4'b0000 ;

endmodule